library verilog;
use verilog.vl_types.all;
entity crc_tb is
end crc_tb;
